library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity shift_direita is
	generic(
		nbits : integer := 4;
		shift : integer := 1
	);
	port(
		op_a, op_b : in std_logic_vector(nbits-1 downto 0);
		resultado : out std_logic_vector(nbits-1 downto 0)
	);
end shift_direita;

architecture comportamento of shift_direita is
begin
	resultado <= std_logic_vector(shift_right(unsigned(op_a), shift));
end comportamento;
